module fa (cout,sum,a,b,c); //6
input a,b,c;
output cout,sum;

ha HA1(c0,s0,a,b);
ha HA2(c1,sum,s0,c);
ha HA3(ignored,cout,c1,c0);

endmodule
